module alu_control_unit(Inp,Out);
input [15:0]Inp;
output [6:0]Out;



assign Out=(Inp[15:12]==4'b1000)?7'b000_0010:
(Inp[15:11]==5'b10011)?7'b000_0100:
(Inp[15:11]==5'b10010)?7'b000_1000:
(Inp[15:11]==5'b10110)?7'b001_0000:
(Inp[15:11]==5'b10101)?7'b010_0000:
(Inp[15:11]==5'b10100)?7'b100_0000:
(Inp[15:14]==2'b0||
Inp[15:14]==2'b01)||
(Inp[15:14]==2'b11&&!(Inp[13:11]==3'b111))?7'b000_0001:7'b0;

endmodule

